module tb;
 initial begin
   $display("Hi dharma welcome,be the truth as much as possible");
  $display("good job man");
 end
endmodule


